
module CPU();
//	input clk
//)
//	wire register_file_A_output
//	
//	
//	
//	
//	FUCKER mem();

endmodule
