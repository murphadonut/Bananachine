module shifter();

endmodule 