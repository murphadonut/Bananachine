
// for branch displacement
// set alu_A_src to 0 for accessing the pc
// set alu_B_src to 1 for immediate value from instruction to add to pc
// set pc_src to 0 for result from alu


// reg B will be used to store stuff to memory
// dont need dual port ram for external memory, just single port will do

module CPU();
//	input clk
//)
//	wire register_file_A_output
//	
//	
//	
//	
//	FUCKER mem();

endmodule
